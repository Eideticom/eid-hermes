`ifndef CONSTANTS
`define CONSTANTS

typedef bit signed [127:0] longlongint;

`endif