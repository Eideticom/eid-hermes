`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Simple module to compute the logical AND of two 32 bit inputs
//////////////////////////////////////////////////////////////////////////////////


module And_32bit(
    input [31:0] a,
    input [31:0] b,
    output [31:0] c
    );
    
    assign c = a&b; 
    
endmodule
